//--------------------------------------------------------------------
//
// Author      : Omkar Girish Kamath
// Date        : April 6th, 2024
// File        : g2b
// Description : gray to binary converter file
//--------------------------------------------------------------------

module g2b (
	    in,
	    out
	    );
   
   //`include "parameter.v"
   //parameter N = $clog2(D);
   parameter N = 9;
   
   //--------------------------------------------------------------------
   // inputs
   //--------------------------------------------------------------------
   input wire [N-1:0] in;
   
   //--------------------------------------------------------------------
   // outputs
   //--------------------------------------------------------------------
   output reg [N-1:0] out;
   
   //--------------------------------------------------------------------
   // internals
   //--------------------------------------------------------------------
   integer 	    i;
   
   //--------------------------------------------------------------------
   // module
   //--------------------------------------------------------------------
   always @(*)
     begin
	out[N-1] = in[N-1];                    // b_(n) = g_(n)
	for (i = N-2; i >= 0; i = i - 1)   
	  out[i] = out[i + 1] ^ in[i];     // b_(i) = b_(i+1) ^ g_(i)
     end
   
endmodule
